module beeper(
input beep,
output bell
);

assign bell = beep;

endmodule
